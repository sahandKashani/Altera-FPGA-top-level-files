-- #############################################################################
-- DE0_Nano_SoC_LT24_top_level.vhd
--
-- BOARD         : DE0-Nano-SoC from Terasic
-- Author        : Sahand Kashani-Akhavan from Terasic documentation
-- Revision      : 1.1
-- Creation date : 11/06/2015
--
-- Syntax Rule : GROUP_NAME_N[bit]
--
-- GROUP : specify a particular interface (ex: SDR_)
-- NAME  : signal name (ex: CONFIG, D, ...)
-- bit   : signal index
-- _N    : to specify an active-low signal
-- #############################################################################

library ieee;
use ieee.std_logic_1164.all;

entity DE0_Nano_SoC_top_level is
    port(
        -- ADC
        ADC_CONVST               : out   std_logic;
        ADC_SCK                  : out   std_logic;
        ADC_SDI                  : out   std_logic;
        ADC_SDO                  : in    std_logic;

        -- ARDUINO
        ARDUINO_IO               : inout std_logic_vector(15 downto 0);
        ARDUINO_RESET_N          : inout std_logic;

        -- CLOCK
        FPGA_CLK1_50             : in    std_logic;
        FPGA_CLK2_50             : in    std_logic;
        FPGA_CLK3_50             : in    std_logic;

        -- KEY
        KEY_N                    : in    std_logic_vector(1 downto 0);

        -- LED
        LED                      : out   std_logic_vector(7 downto 0);

        -- SW
        SW                       : in    std_logic_vector(3 downto 0);

        -- GPIO_0
        GPIO_0_LT24_ADC_BUSY     : in    std_logic;
        GPIO_0_LT24_ADC_CS_N     : out   std_logic;
        GPIO_0_LT24_ADC_DCLK     : out   std_logic;
        GPIO_0_LT24_ADC_DIN      : out   std_logic;
        GPIO_0_LT24_ADC_DOUT     : in    std_logic;
        GPIO_0_LT24_ADC_PENIRQ_N : in    std_logic;
        GPIO_0_LT24_CS_N         : out   std_logic;
        GPIO_0_LT24_D            : out   std_logic_vector(15 downto 0);
        GPIO_0_LT24_LCD_ON       : out   std_logic;
        GPIO_0_LT24_RD_N         : out   std_logic;
        GPIO_0_LT24_RESET_N      : out   std_logic;
        GPIO_0_LT24_RS           : out   std_logic;
        GPIO_0_LT24_WR_N         : out   std_logic;

        -- GPIO_1
        GPIO_1                   : inout std_logic_vector(35 downto 0);

        -- HPS
        HPS_CONV_USB_N           : inout std_logic;
        HPS_DDR3_ADDR            : out   std_logic_vector(14 downto 0);
        HPS_DDR3_BA              : out   std_logic_vector(2 downto 0);
        HPS_DDR3_CAS_N           : out   std_logic;
        HPS_DDR3_CK_N            : out   std_logic;
        HPS_DDR3_CK_P            : out   std_logic;
        HPS_DDR3_CKE             : out   std_logic;
        HPS_DDR3_CS_N            : out   std_logic;
        HPS_DDR3_DM              : out   std_logic_vector(3 downto 0);
        HPS_DDR3_DQ              : inout std_logic_vector(31 downto 0);
        HPS_DDR3_DQS_N           : inout std_logic_vector(3 downto 0);
        HPS_DDR3_DQS_P           : inout std_logic_vector(3 downto 0);
        HPS_DDR3_ODT             : out   std_logic;
        HPS_DDR3_RAS_N           : out   std_logic;
        HPS_DDR3_RESET_N         : out   std_logic;
        HPS_DDR3_RZQ             : in    std_logic;
        HPS_DDR3_WE_N            : out   std_logic;
        HPS_ENET_GTX_CLK         : out   std_logic;
        HPS_ENET_INT_N           : inout std_logic;
        HPS_ENET_MDC             : out   std_logic;
        HPS_ENET_MDIO            : inout std_logic;
        HPS_ENET_RX_CLK          : in    std_logic;
        HPS_ENET_RX_DATA         : in    std_logic_vector(3 downto 0);
        HPS_ENET_RX_DV           : in    std_logic;
        HPS_ENET_TX_DATA         : out   std_logic_vector(3 downto 0);
        HPS_ENET_TX_EN           : out   std_logic;
        HPS_GSENSOR_INT          : inout std_logic;
        HPS_I2C0_SCLK            : inout std_logic;
        HPS_I2C0_SDAT            : inout std_logic;
        HPS_I2C1_SCLK            : inout std_logic;
        HPS_I2C1_SDAT            : inout std_logic;
        HPS_KEY_N                : inout std_logic;
        HPS_LED                  : inout std_logic;
        HPS_LTC_GPIO             : inout std_logic;
        HPS_SD_CLK               : out   std_logic;
        HPS_SD_CMD               : inout std_logic;
        HPS_SD_DATA              : inout std_logic_vector(3 downto 0);
        HPS_SPIM_CLK             : out   std_logic;
        HPS_SPIM_MISO            : in    std_logic;
        HPS_SPIM_MOSI            : out   std_logic;
        HPS_SPIM_SS              : inout std_logic;
        HPS_UART_RX              : in    std_logic;
        HPS_UART_TX              : out   std_logic;
        HPS_USB_CLKOUT           : in    std_logic;
        HPS_USB_DATA             : inout std_logic_vector(7 downto 0);
        HPS_USB_DIR              : in    std_logic;
        HPS_USB_NXT              : in    std_logic;
        HPS_USB_STP              : out   std_logic
    );
end entity DE0_Nano_SoC_top_level;

architecture rtl of DE0_Nano_SoC_top_level is

begin

end;
